library verilog;
use verilog.vl_types.all;
entity FPU_tb is
end FPU_tb;
